`timescale 1ns / 1ps
/*********************************************************
 * File Name: MIPS_top.v
 * Project: MIPS ISA Processor - Senior Project
 * Designer: Steven Sallack & Michael Diep
 * Email: Steven.Sallack@gmail.com // michaelkhangdiep@gmail.com
 * Rev. Date: 4/23/2018
 *
 * Purpose: This module instantiates the necessary modules needed to
 *          have a working pipelined MIPS processor. The interrupt
 *          is serviced by saving the PC to $31 and
 *          retrieving the ISR location from memory. When the ISR is 
 *          finished and a JR instruction is reached, it loads the PC
 *          with the contents of $31 and resumes fetching and executing 
 *          instructions.
 *                 
 *          Data memory bus should be connected to D_out input. 
 *          I/O data bus should be connected to the IO_IN input;
 *
 * Notes: Rev. 3/21/18  - updated header and adjusted comments
 *        
 *        Rev. 4/21/18  - implemented modules 1-13 and updated header
 *********************************************************/
module MIPS_top(clk, rst, intr, D_out, IO_IN, 
                inta, EX_MEM, RTOUT, ALU_OUT, EX_MEM_IO_SEL);
input clk, rst, intr;
input [31:0] D_out, IO_IN;
output inta;
output [49:0] EX_MEM; 
output [31:0] RTOUT, ALU_OUT;
output [2:0] EX_MEM_IO_SEL;

//wire interconnections
wire [31:0] IR_out, PC_out, SE_16, ALU_OUT, D_in, D_out, PC_in, 
            DY, D_OUT, MEM2REG, RTOUT, RSB, RTB, RFD, JR_RS, IO_IN, TO_PC_IN;

//control signal from PMCU
wire int_ack;
wire [1:0]  m2r;
wire D_en, HILO_ld, T_sel;
wire [1:0] D_sel;
wire [2:0] Y_sel, RFD_sel;
wire [4:0] FS;
wire dm_cs, dm_rd, dm_wr;

wire [17:0] CONTROL;

wire [1:0] ForwardA, ForwardB;

wire [1:0] PC_SEL;

wire ifjump, ifjr, dojr, doBranch;

wire [4:0] TO_EX_MEM_DEST; // rt if I type, rd if R type
wire IloRhi; //I or R type instruction
wire Break; //generated to end the simulation
wire SW_HI, OUT_HI; 
wire isBranch, stall, io_cs, io_rd, io_wr, INT_INPROG;

wire ns_N, ns_Z, ns_C, ns_V, ns_IE;

//registers
reg ps_N, ps_Z, ps_C, ps_V, ps_IE;
reg [49:0] ID_EX, EX_MEM, MEM_WB; //pipeline registers
reg [31:0] MEM_WB_ALU_OUT, MEM_OUT, IO_MEM_OUT, RT_MEM, ID_EX_SE_16;
reg [31:0] IF_ID_PC, ID_EX_PC, EX_MEM_PC, MEM_WB_PC; //pipeline registers for PC
reg [2:0] ID_EX_RFD, EX_MEM_RFD, MEM_WB_RFD, ID_EX_IO_SEL, EX_MEM_IO_SEL;
reg [4:0] EX_MEM_DEST, MEM_WB_DEST; //dest reg of inst-1 and inst-2
reg       ID_EX_INTR, EX_MEM_INTR, MEM_WB_INTR;



   // synchronous flags register assignment
   always @ (posedge clk or posedge rst)
      if (rst)
         {ps_N,ps_Z,ps_C, ps_V, ps_IE} <= 5'b0;
      else
         {ps_N,ps_Z,ps_C, ps_V, ps_IE} <= {ns_N,ns_Z,ns_C,ns_V,ns_IE};
         
    //pipeline registers contain full instruction and 
    //   control signals generated by Pipelined_MCU
    //IR_out is first stage of pipeline registers       
   always @(posedge clk or posedge rst)
      if (rst)
         {ID_EX, EX_MEM, MEM_WB} <= 150'h0; else 
      if (stall) {ID_EX, EX_MEM, MEM_WB} <= {50'h0, ID_EX, EX_MEM}; else
      if (intr & ps_IE)  {ID_EX, EX_MEM, MEM_WB} <= 
                         {{32'b0,18'b01_0110_0001_0101_0101}, ID_EX, EX_MEM}; else
         {ID_EX, EX_MEM, MEM_WB} <= {{IR_out,CONTROL}, ID_EX, EX_MEM};
      
         //pipeline registers for PC
   always @(posedge clk or posedge rst)
      if (rst)
      {IF_ID_PC, ID_EX_PC, EX_MEM_PC, MEM_WB_PC} <= 128'h0; else
      {IF_ID_PC, ID_EX_PC, EX_MEM_PC, MEM_WB_PC} <= 
                                    {PC_out, IF_ID_PC, ID_EX_PC, EX_MEM_PC};
    
      //ALU_OUT buffer register for WB
   always @(posedge clk or posedge rst) 
      if (rst) 
            MEM_WB_ALU_OUT <= 32'h0; else
            MEM_WB_ALU_OUT <= ALU_OUT;
       
         //MEM output register for WB
    always @(posedge clk or posedge rst)
      if (rst) 
            {MEM_OUT, IO_MEM_OUT} <= 64'h0; else
            {MEM_OUT, IO_MEM_OUT} <= {D_out, IO_IN};
    
    //reg for IO control signals
    always @(posedge clk or posedge rst)
      if (rst)
         {ID_EX_IO_SEL, EX_MEM_IO_SEL} <= 6'b0; else
         {ID_EX_IO_SEL, EX_MEM_IO_SEL} <= 
                     {{io_cs, io_wr, io_rd}, ID_EX_IO_SEL};
    
     //pipe reg's for RFD_sel 
     always @(posedge clk or posedge rst)
      if (rst) {ID_EX_RFD, EX_MEM_RFD, MEM_WB_RFD} <= 9'h0; else if
         (intr & ps_IE){ID_EX_RFD, EX_MEM_RFD, MEM_WB_RFD} <= 
                                 {3'h3, ID_EX_RFD, EX_MEM_RFD}; else
               {ID_EX_RFD, EX_MEM_RFD, MEM_WB_RFD} <= 
                                 {RFD_sel, ID_EX_RFD, EX_MEM_RFD};
               
     //pipe reg's for interrupt signals
     always @(posedge clk or posedge rst)
      if (rst) 
               {ID_EX_INTR, EX_MEM_INTR, MEM_WB_INTR} <= 3'h0;
          else if (ps_IE) 
               {ID_EX_INTR, EX_MEM_INTR, MEM_WB_INTR} <= 
                                          {intr, ID_EX_INTR, EX_MEM_INTR};
       
     //pipe reg's for destination registers
     always @(posedge clk or posedge rst)
      if (rst) 
      {EX_MEM_DEST, MEM_WB_DEST} <= 10'h0; else
      if (SW_HI | OUT_HI) //need to make store word / output put 0s
      {EX_MEM_DEST, MEM_WB_DEST} <= {5'h0, EX_MEM_DEST}; else 
      {EX_MEM_DEST, MEM_WB_DEST} <= {TO_EX_MEM_DEST, EX_MEM_DEST};  
       
     //pipeline the sign extension
     always @(posedge clk or posedge rst)
      if (rst) ID_EX_SE_16 <= 32'b0; else
               ID_EX_SE_16 <= SE_16;
               
       //destination register for forwarding, rt if i type, rd if r type
    assign TO_EX_MEM_DEST = (ID_EX[49:44] == 0)? ID_EX[33:29] : //R-Type - pass Rd
                            (ID_EX[49:44] != 0)? ID_EX[38:34] : //I-Type - pass Rt               
                                                  5'h0; //default (j type)
                                                  
     //determine if instruction about to be executed is R or I type
    assign IloRhi = (ID_EX[49:44] == 6'h0);
     //determine if instruction about to be executed is a SW
    assign SW_HI  = (ID_EX[49:44] == 6'h2B);
    //determine if instruction about to be executed is an output
    assign OUT_HI = (ID_EX[49:44] == 6'h1D);
    
    //need stall for LW->SW (stall if next instruction uses destination of LW)
    assign stall = (ID_EX[14] & ((ID_EX[38:34] == IR_out[25:21]) 
                     | (ID_EX[38:34] == IR_out[20:16])));
     
     //control net determined in decode
    assign CONTROL = {m2r,dm_wr,dm_rd,dm_cs,Y_sel,HILO_ld,FS,T_sel,D_sel,D_en};
    
    //ALU_OUT, memory output, or IO output data
    assign MEM2REG = (MEM_WB[17:16] == 2'b00) ? MEM_WB_ALU_OUT : 
                     (MEM_WB[17:16] == 2'b01) ? MEM_OUT :      
                     (MEM_WB[17:16] == 2'b10) ? IO_MEM_OUT : MEM_WB_ALU_OUT; 
    
    assign ifjump = ((IR_out[31:26] == 6'h02) 
                  | (IR_out[31:26] == 6'h03)); //is a jump or jal
                  
    assign dojr = ((ID_EX[49:44]==6'h0) 
                  & (ID_EX[23:18] == 6'h08)); //is a jr
                  
    assign ifjr = ((IR_out[31:26]==6'h0) 
                  & (IR_out[5:0] == 6'h08)); //see a jr
    
    //dont inc the pc
    assign NO_INC = (ifjump | doBranch | ifjr | dojr 
                     | isBranch | stall | INT_INPROG); 
    
    //used to save PC from a pipeline PC register
    assign RFD = (MEM_WB_RFD == 3'h0)? MEM2REG : 
                 (MEM_WB_RFD == 3'h1)? IF_ID_PC:
                 (MEM_WB_RFD == 3'h2)? ID_EX_PC:
                 (MEM_WB_RFD == 3'h3)? EX_MEM_PC:
                 (MEM_WB_RFD == 3'h4)? MEM_WB_PC:
                                    MEM2REG;
    
    //assigned if is jump or jr (branch uses default 0)
    assign PC_SEL = ({ifjump, dojr, MEM_WB_INTR} == 3'b000)? 2'b00 :
                    ({ifjump, dojr, MEM_WB_INTR} == 3'b010)? 2'b10 :
                    ({ifjump, dojr, MEM_WB_INTR} == 3'b100)? 2'b01 :
                    ({ifjump, dojr, MEM_WB_INTR} == 3'b100)? 2'b00 :
                    ({ifjump, dojr, MEM_WB_INTR} == 3'b001)? 2'b10 : 2'b00;
    
    //if the interrupt is being serviced
    assign INT_INPROG = (ps_IE & (intr | ID_EX_INTR | EX_MEM_INTR | MEM_WB_INTR));
    
    //need to take RSB to PC for JR, else using MEM2REG
    assign TO_PC_IN = (dojr)? RSB : MEM2REG; 
    
    //acknowledge the interrupt 
    assign inta = (MEM_WB_INTR);
    
   BreakCounter BreakC (
      .clk(clk),
      .rst(rst),
      .IR(IR_out[31:0]),
      .done(Break)
      );
      
   ForwardingUnit FU (
      .isBranch(isBranch),
      .IloRhi(IloRhi),
      .OUT_HI(OUT_HI),
      .SW_HI(SW_HI),
      .RS(ID_EX[43:39]),
      .RT(ID_EX[38:34]),
      .RD_M1(EX_MEM_DEST),
      .RD_M2(MEM_WB_DEST),
      .FA(ForwardA),
      .FB(ForwardB)
      );
                          
	Instruction_Unit IU (
		.clk(clk), 
		.rst(rst), 
		.im_cs(1'b1), 
		.im_wr(1'b0), 
		.im_rd(1'b1), 
		.pc_sel(PC_SEL), 
		.pc_ld((ifjump | doBranch | dojr | (ps_IE & MEM_WB_INTR))), 
		.pc_inc(~NO_INC), 
		.ir_ld(~(ifjump | doBranch | isBranch | stall | ifjr | dojr | INT_INPROG)), 
		.PC_in(TO_PC_IN), 
		.PC_out(PC_out), 
		.IR_out(IR_out), 
		.SE_16(SE_16),
      .RSB(JR_RS), 
      .nop(ifjump | doBranch | isBranch | ifjr), 
      .ID_EX_SE_16(ID_EX_SE_16)     
	);
   
   BranchControl BC (
         .IRF(IR_out),
         .IREX(ID_EX[49:18]),
         .RS(RSB), 
         .RT(RTB), 
         .doBranch(doBranch),
         .isBranch(isBranch)
         );

	Integer_Datapath IDP (
		.clk(clk),
      .rst(rst),
      .RSB(RSB), 
      .RTB(RTB), 
      .RTOUT(RTOUT), 
      .D(RFD), 
      .FS(ID_EX[8:4]),
      .shamt(ID_EX[28:24]),
      .S_addr(IR_out[25:21]),
      .T_addr(IR_out[20:16]),
      .D_addr0(MEM_WB[33:29]), //$rd
      .D_addr1(MEM_WB[38:34]),  //$rt
      .D_en(MEM_WB[0]),
      .DT(ID_EX_SE_16),
      .HILO_ld(ID_EX[9]),
      .T_sel(ID_EX[3]),
      .DY(D_out),
      .PC_in(IR_out),
      .Y_sel(EX_MEM[12:10]),
      .D_sel(MEM_WB[2:1]), 
		.ALU_OUT(ALU_OUT), 
		.C(ns_C), 
		.V(ns_V), 
		.N(ns_N), 
		.Z(ns_Z),
      .FWDA_SEL(ForwardA),
      .FWDB_SEL(ForwardB),
      .EX_MEM_FWD(ALU_OUT),
      .MEM_WB_FWD(MEM2REG),
      .RFS2RS(JR_RS),
      .IO_IN(IO_IN)
	);  
          
   	Pipelined_MCU PMCU(
		.intr(intr), 
      .IE(ps_IE),
		.IR(IR_out), 
      .FS(FS),
		.D_en(D_en), 
		.D_sel(D_sel), 
		.T_sel(T_sel), 
		.HILO_ld(HILO_ld), 
		.Y_sel(Y_sel), 
		.dm_cs(dm_cs), 
		.dm_rd(dm_rd), 
		.dm_wr(dm_wr),
      .new_IE(ns_IE),
      .m2r(m2r),
      .RFD_sel(RFD_sel),
      .io_cs(io_cs),
      .io_wr(io_wr),
      .io_rd(io_rd)
	);

endmodule
